library work;
use work.my_components.all;

